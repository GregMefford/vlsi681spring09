module ALU(A, B, CONTROL, CC, Z, OF);

    input  [15:0] A;       // port A
    input  [15:0] B;       // port B
    input  [ 2:0] CONTROL; // control for ALU
    output [ 2:0] CC;      // pos, neg, zero flags
    output [15:0] Z;       // result
    output        OF;      // overflow
    wire   [16:0] result;  // ALU result


    assign result = alu_out(A, B, CONTROL);
    assign Z = result[15:0];
    assign OF  = result[16];
    assign CC = flags(result);

     function [16:0] alu_out;
           input  [15:0] A,B;
           input  [2:0] CONTROL;
           case (CONTROL)
                   3'b000: alu_out=A+B;              // Add A,B
                   3'b001: alu_out=A&B;              // And A,B
                   3'b010: alu_out=~A;               // Not A
                   3'b100: alu_out=A[7:0] * B[7:0];  // Mul A,B
                   3'b110: alu_out={A[14:0],1'b0};   // Shift Left
                   3'b101: alu_out={A[15],A[15:1]};  // Shift Right (sign extend)
                 default: begin
                             alu_out=17'bX;
                       end    
             endcase  /* {...,...,...} is for the concatenation.
                         {ADD_WITH_CARRY,SUB_WITH_BORROW}==2'b11 is used
                         to force the CARRY==1 for the increment operation */  
       endfunction // end of function "result"

      function [2:0] flags;        // output [pos,neg,zero] flags
          input [16:0] x;
          
            begin

            //initialize flags to zero
            flags[0] = 0;
            flags[1] = 0;
            flags[2] = 0;
            
            // zero flag check for x
            if( x == 0)
            begin
                flags[0] = 1;
            end
            else
            begin
                if(x[16] == 1)
                begin
                    flags[1] = 1;
                    flags[2] = 0;
                end
                else
                begin
                    flags[1] = 0;
                    flags[2] = 1;
                end
            end
            end
      endfunction // end of function "flags"
endmodule
