module RAM_instruction(CLK, ADDRESS, INSTRUCTION);
	input              CLK;
	input      [15: 0] ADDRESS;
	output reg [15: 0] INSTRUCTION;
	
endmodule
