library verilog;
use verilog.vl_types.all;
entity altmult_accum is
    generic(
        width_a         : integer := 2;
        width_b         : integer := 2;
        width_result    : integer := 5;
        input_reg_a     : string  := "CLOCK0";
        input_aclr_a    : string  := "ACLR3";
        input_reg_b     : string  := "CLOCK0";
        input_aclr_b    : string  := "ACLR3";
        port_addnsub    : string  := "PORT_CONNECTIVITY";
        addnsub_reg     : string  := "CLOCK0";
        addnsub_aclr    : string  := "ACLR3";
        addnsub_pipeline_reg: string  := "CLOCK0";
        addnsub_pipeline_aclr: string  := "ACLR3";
        accum_direction : string  := "ADD";
        accum_sload_reg : string  := "CLOCK0";
        accum_sload_aclr: string  := "ACLR3";
        accum_sload_pipeline_reg: string  := "CLOCK0";
        accum_sload_pipeline_aclr: string  := "ACLR3";
        representation_a: string  := "UNSIGNED";
        port_signa      : string  := "PORT_CONNECTIVITY";
        sign_reg_a      : string  := "CLOCK0";
        sign_aclr_a     : string  := "ACLR3";
        sign_pipeline_reg_a: string  := "CLOCK0";
        sign_pipeline_aclr_a: string  := "ACLR3";
        port_signb      : string  := "PORT_CONNECTIVITY";
        representation_b: string  := "UNSIGNED";
        sign_reg_b      : string  := "CLOCK0";
        sign_aclr_b     : string  := "ACLR3";
        sign_pipeline_reg_b: string  := "CLOCK0";
        sign_pipeline_aclr_b: string  := "ACLR3";
        multiplier_reg  : string  := "CLOCK0";
        multiplier_aclr : string  := "ACLR3";
        output_reg      : string  := "CLOCK0";
        output_aclr     : string  := "ACLR3";
        lpm_type        : string  := "altmult_accum";
        lpm_hint        : string  := "UNUSED";
        extra_multiplier_latency: integer := 0;
        extra_accumulator_latency: integer := 0;
        dedicated_multiplier_circuitry: string  := "AUTO";
        dsp_block_balancing: string  := "AUTO";
        intended_device_family: string  := "Stratix";
        accum_round_aclr: string  := "ACLR3";
        accum_round_pipeline_aclr: string  := "ACLR3";
        accum_round_pipeline_reg: string  := "CLOCK0";
        accum_round_reg : string  := "CLOCK0";
        accum_saturation_aclr: string  := "ACLR3";
        accum_saturation_pipeline_aclr: string  := "ACLR3";
        accum_saturation_pipeline_reg: string  := "CLOCK0";
        accum_saturation_reg: string  := "CLOCK0";
        accum_sload_upper_data_aclr: string  := "ACLR3";
        accum_sload_upper_data_pipeline_aclr: string  := "ACLR3";
        accum_sload_upper_data_pipeline_reg: string  := "CLOCK0";
        accum_sload_upper_data_reg: string  := "CLOCK0";
        mult_round_aclr : string  := "ACLR3";
        mult_round_reg  : string  := "CLOCK0";
        mult_saturation_aclr: string  := "ACLR3";
        mult_saturation_reg: string  := "CLOCK0";
        input_source_a  : string  := "DATAA";
        input_source_b  : string  := "DATAB";
        width_upper_data: integer := 1;
        multiplier_rounding: string  := "NO";
        multiplier_saturation: string  := "NO";
        accumulator_rounding: string  := "NO";
        accumulator_saturation: string  := "NO";
        port_mult_is_saturated: string  := "UNUSED";
        port_accum_is_saturated: string  := "UNUSED"
    );
    port(
        dataa           : in     vl_logic_vector;
        datab           : in     vl_logic_vector;
        scanina         : in     vl_logic_vector;
        scaninb         : in     vl_logic_vector;
        sourcea         : in     vl_logic;
        sourceb         : in     vl_logic;
        accum_sload_upper_data: in     vl_logic_vector;
        addnsub         : in     vl_logic;
        accum_sload     : in     vl_logic;
        signa           : in     vl_logic;
        signb           : in     vl_logic;
        clock0          : in     vl_logic;
        clock1          : in     vl_logic;
        clock2          : in     vl_logic;
        clock3          : in     vl_logic;
        ena0            : in     vl_logic;
        ena1            : in     vl_logic;
        ena2            : in     vl_logic;
        ena3            : in     vl_logic;
        aclr0           : in     vl_logic;
        aclr1           : in     vl_logic;
        aclr2           : in     vl_logic;
        aclr3           : in     vl_logic;
        result          : out    vl_logic_vector;
        overflow        : out    vl_logic;
        scanouta        : out    vl_logic_vector;
        scanoutb        : out    vl_logic_vector;
        mult_round      : in     vl_logic;
        mult_saturation : in     vl_logic;
        accum_round     : in     vl_logic;
        accum_saturation: in     vl_logic;
        mult_is_saturated: out    vl_logic;
        accum_is_saturated: out    vl_logic
    );
end altmult_accum;
