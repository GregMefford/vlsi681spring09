module Execution(
	input	[2:0]  ALU_CONTROL,
	input	       ALU_MuxA,
	input	[2:0]  ALU_MuxB,
	input	[15:0] PC,
	input	[15:0] IR,
	input	[15:0] RS1_DATA,
	input	[15:0] RS2_DATA,
	output	       N,
	output	       Z,
	output	       P,
	output         OF,
	output	[15:0] Y
);

wire	[15:0] IMM5_SE;
wire	[15:0] ALU_A;
wire	[15:0] ALU_B;
wire    [ 2:0] NPZ;

assign ALU_A = (ALU_MuxA) ? RS1_DATA : PC;
assign N = NPZ[2];
assign P = NPZ[1];
assign Z = NPZ[0];

assign ALU_B = alu_muxb(IR, RS2_DATA, ALU_MuxB);
function [15:0] alu_muxb;
	input [15:0] IR;
	input [15:0] RS2_DATA;
	input [ 2:0] ALU_MuxB;
	if(ALU_MuxB[2]) begin
	  case(ALU_MuxB[1:0])
	    'b00: alu_muxb = {{11{IR[ 4]}}, IR[ 4:0]}; // IMM5
	    'b01: alu_muxb = {{10{IR[ 5]}}, IR[ 5:0]}; // Offset6
	    'b10: alu_muxb = {{ 7{IR[ 8]}}, IR[ 8:0]}; // Offset9
	    'b11: alu_muxb = {{ 5{IR[10]}}, IR[10:0]}; // Offset11
	    default: alu_muxb = 16'bX;
	  endcase
	end
	else alu_muxb = RS2_DATA;
endfunction // alu_muxb

ALU	ALU_inst(
	.A(ALU_A),
	.B(ALU_B),
	.CONTROL(ALU_CONTROL),

  .OF(OF),
	.CC(NPZ),
	.Z(Y)
);

endmodule
