library verilog;
use verilog.vl_types.all;
entity altdq_dqs is
    generic(
        delay_buffer_mode: string  := "LOW";
        delay_dqs_enable_by_half_cycle: string  := "FALSE";
        intended_device_family: string  := "UNUSED";
        dq_half_rate_use_dataoutbypass: string  := "FALSE";
        dq_input_reg_async_mode: string  := "NONE";
        dq_input_reg_clk_source: string  := "DQS_BUS";
        dq_input_reg_mode: string  := "NONE";
        dq_input_reg_power_up: string  := "LOW";
        dq_input_reg_sync_mode: string  := "NONE";
        dq_input_reg_use_clkn: string  := "FALSE";
        dq_ipa_add_input_cycle_delay: string  := "FALSE";
        dq_ipa_add_phase_transfer_reg: string  := "FALSE";
        dq_ipa_bypass_output_register: string  := "FALSE";
        dq_ipa_invert_phase: string  := "FALSE";
        dq_ipa_phase_setting: integer := 0;
        dq_oe_reg_async_mode: string  := "NONE";
        dq_oe_reg_mode  : string  := "NONE";
        dq_oe_reg_power_up: string  := "LOW";
        dq_oe_reg_sync_mode: string  := "NONE";
        dq_output_reg_async_mode: string  := "NONE";
        dq_output_reg_mode: string  := "NONE";
        dq_output_reg_power_up: string  := "LOW";
        dq_output_reg_sync_mode: string  := "NONE";
        dqs_ctrl_latches_enable: string  := "FALSE";
        dqs_delay_chain_delayctrlin_source: string  := "CORE";
        dqs_delay_chain_phase_setting: integer := 0;
        dqs_dqsn_mode   : string  := "NONE";
        dqs_enable_ctrl_add_phase_transfer_reg: string  := "FALSE";
        dqs_enable_ctrl_invert_phase: string  := "FALSE";
        dqs_enable_ctrl_phase_setting: integer := 0;
        dqs_input_frequency: string  := "UNUSED";
        dqs_oe_reg_async_mode: string  := "NONE";
        dqs_oe_reg_mode : string  := "NONE";
        dqs_oe_reg_power_up: string  := "LOW";
        dqs_oe_reg_sync_mode: string  := "NONE";
        dqs_offsetctrl_enable: string  := "FALSE";
        dqs_output_reg_async_mode: string  := "NONE";
        dqs_output_reg_mode: string  := "NONE";
        dqs_output_reg_power_up: string  := "LOW";
        dqs_output_reg_sync_mode: string  := "NONE";
        dqs_phase_shift : integer := 0;
        io_clock_divider_clk_source: string  := "CORE";
        io_clock_divider_invert_phase: string  := "FALSE";
        io_clock_divider_phase_setting: integer := 0;
        level_dqs_enable: string  := "FALSE";
        number_of_bidir_dq: integer := 1;
        number_of_clk_divider: integer := 1;
        number_of_input_dq: integer := 1;
        number_of_output_dq: integer := 1;
        oct_reg_mode    : string  := "NONE";
        use_dq_input_delay_chain: string  := "FALSE";
        use_dq_ipa      : string  := "FALSE";
        use_dq_ipa_phasectrlin: string  := "TRUE";
        use_dq_oe_delay_chain1: string  := "FALSE";
        use_dq_oe_delay_chain2: string  := "FALSE";
        use_dq_oe_path  : string  := "FALSE";
        use_dq_output_delay_chain1: string  := "FALSE";
        use_dq_output_delay_chain2: string  := "FALSE";
        use_dqs         : string  := "FALSE";
        use_dqs_delay_chain: string  := "FALSE";
        use_dqs_delay_chain_phasectrlin: string  := "FALSE";
        use_dqs_enable  : string  := "FALSE";
        use_dqs_enable_ctrl: string  := "FALSE";
        use_dqs_enable_ctrl_phasectrlin: string  := "TRUE";
        use_dqs_input_delay_chain: string  := "FALSE";
        use_dqs_input_path: string  := "FALSE";
        use_dqs_oe_delay_chain1: string  := "FALSE";
        use_dqs_oe_delay_chain2: string  := "FALSE";
        use_dqs_oe_path : string  := "FALSE";
        use_dqs_output_delay_chain1: string  := "FALSE";
        use_dqs_output_delay_chain2: string  := "FALSE";
        use_dqs_output_path: string  := "FALSE";
        use_dqsbusout_delay_chain: string  := "FALSE";
        use_dqsenable_delay_chain: string  := "FALSE";
        use_dynamic_oct : string  := "FALSE";
        use_half_rate   : string  := "FALSE";
        use_io_clock_divider_masterin: string  := "FALSE";
        use_io_clock_divider_phasectrlin: string  := "TRUE";
        use_oct_delay_chain1: string  := "FALSE";
        use_oct_delay_chain2: string  := "FALSE";
        lpm_hint        : string  := "UNUSED";
        lpm_type        : string  := "altdq_dqs"
    );
    port(
        bidir_dq_areset : in     vl_logic_vector;
        bidir_dq_hr_oct_in: in     vl_logic_vector;
        bidir_dq_hr_oe_in: in     vl_logic_vector;
        bidir_dq_hr_output_data_in: in     vl_logic_vector;
        bidir_dq_input_data_in: in     vl_logic_vector;
        bidir_dq_io_config_ena: in     vl_logic_vector;
        bidir_dq_oct_in : in     vl_logic_vector;
        bidir_dq_oe_in  : in     vl_logic_vector;
        bidir_dq_output_data_in: in     vl_logic_vector;
        bidir_dq_output_data_in_high: in     vl_logic_vector;
        bidir_dq_output_data_in_low: in     vl_logic_vector;
        bidir_dq_sreset : in     vl_logic_vector;
        config_clk      : in     vl_logic;
        config_datain   : in     vl_logic;
        config_update   : in     vl_logic;
        core_delayctrlin: in     vl_logic_vector(5 downto 0);
        dll_delayctrlin : in     vl_logic_vector(5 downto 0);
        dq_hr_output_reg_clk: in     vl_logic;
        dq_input_reg_clk: in     vl_logic;
        dq_input_reg_clkena: in     vl_logic;
        dq_ipa_clk      : in     vl_logic;
        dq_output_reg_clk: in     vl_logic;
        dq_output_reg_clkena: in     vl_logic;
        dqs_areset      : in     vl_logic;
        dqs_config_ena  : in     vl_logic;
        dqs_enable_ctrl_clk: in     vl_logic;
        dqs_enable_ctrl_hr_datainhi: in     vl_logic;
        dqs_enable_ctrl_hr_datainlo: in     vl_logic;
        dqs_enable_ctrl_in: in     vl_logic;
        dqs_enable_in   : in     vl_logic;
        dqs_hr_oct_in   : in     vl_logic_vector(1 downto 0);
        dqs_hr_oe_in    : in     vl_logic_vector(1 downto 0);
        dqs_hr_output_data_in: in     vl_logic_vector(3 downto 0);
        dqs_hr_output_reg_clk: in     vl_logic;
        dqs_input_data_in: in     vl_logic;
        dqs_io_config_ena: in     vl_logic;
        dqs_oct_in      : in     vl_logic;
        dqs_oe_in       : in     vl_logic;
        dqs_output_data_in: in     vl_logic;
        dqs_output_data_in_high: in     vl_logic;
        dqs_output_data_in_low: in     vl_logic;
        dqs_output_reg_clk: in     vl_logic;
        dqs_output_reg_clkena: in     vl_logic;
        dqs_sreset      : in     vl_logic;
        dqsn_areset     : in     vl_logic;
        dqsn_hr_oct_in  : in     vl_logic_vector(1 downto 0);
        dqsn_hr_oe_in   : in     vl_logic_vector(1 downto 0);
        dqsn_hr_output_data_in: in     vl_logic_vector(3 downto 0);
        dqsn_input_data_in: in     vl_logic;
        dqsn_io_config_ena: in     vl_logic;
        dqsn_oct_in     : in     vl_logic;
        dqsn_oe_in      : in     vl_logic;
        dqsn_output_data_in: in     vl_logic;
        dqsn_output_data_in_high: in     vl_logic;
        dqsn_output_data_in_low: in     vl_logic;
        dqsn_sreset     : in     vl_logic;
        dqsupdateen     : in     vl_logic;
        hr_oct_reg_clk  : in     vl_logic;
        input_dq_areset : in     vl_logic_vector;
        input_dq_hr_oct_in: in     vl_logic_vector;
        input_dq_input_data_in: in     vl_logic_vector;
        input_dq_io_config_ena: in     vl_logic_vector;
        input_dq_oct_in : in     vl_logic_vector;
        input_dq_sreset : in     vl_logic_vector;
        io_clock_divider_clk: in     vl_logic;
        io_clock_divider_masterin: in     vl_logic;
        oct_reg_clk     : in     vl_logic;
        offsetctrlin    : in     vl_logic_vector(5 downto 0);
        output_dq_areset: in     vl_logic_vector;
        output_dq_hr_oct_in: in     vl_logic_vector;
        output_dq_hr_oe_in: in     vl_logic_vector;
        output_dq_hr_output_data_in: in     vl_logic_vector;
        output_dq_io_config_ena: in     vl_logic_vector;
        output_dq_oct_in: in     vl_logic_vector;
        output_dq_oe_in : in     vl_logic_vector;
        output_dq_output_data_in: in     vl_logic_vector;
        output_dq_output_data_in_high: in     vl_logic_vector;
        output_dq_output_data_in_low: in     vl_logic_vector;
        output_dq_sreset: in     vl_logic_vector;
        bidir_dq_hr_input_data_out: out    vl_logic_vector;
        bidir_dq_input_data_out: out    vl_logic_vector;
        bidir_dq_input_data_out_high: out    vl_logic_vector;
        bidir_dq_input_data_out_low: out    vl_logic_vector;
        bidir_dq_oct_out: out    vl_logic_vector;
        bidir_dq_oe_out : out    vl_logic_vector;
        bidir_dq_output_data_out: out    vl_logic_vector;
        dqs_bus_out     : out    vl_logic;
        dqs_input_data_out: out    vl_logic;
        dqs_oct_out     : out    vl_logic;
        dqs_oe_out      : out    vl_logic;
        dqs_output_data_out: out    vl_logic;
        dqsn_bus_out    : out    vl_logic;
        dqsn_input_data_out: out    vl_logic;
        dqsn_oct_out    : out    vl_logic;
        dqsn_oe_out     : out    vl_logic;
        dqsn_output_data_out: out    vl_logic;
        input_dq_hr_input_data_out: out    vl_logic_vector;
        input_dq_input_data_out: out    vl_logic_vector;
        input_dq_input_data_out_high: out    vl_logic_vector;
        input_dq_input_data_out_low: out    vl_logic_vector;
        input_dq_oct_out: out    vl_logic_vector;
        io_clock_divider_clkout: out    vl_logic_vector;
        io_clock_divider_slaveout: out    vl_logic;
        output_dq_oct_out: out    vl_logic_vector;
        output_dq_oe_out: out    vl_logic_vector;
        output_dq_output_data_out: out    vl_logic_vector
    );
end altdq_dqs;
